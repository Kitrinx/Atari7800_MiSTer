-------------------------------------------------------------------------------
--
--   Copyright (C) 2005
--
--   Title     :  Atari 2600 TIA control logic and playfield generation
--
--   Author    :  Ed Henciak 
--
--   Notes     :  This component ties together everything for
--                horizontal sync control, playfield logic, and 
--                motion control.  This logic basically controls
--                clocking of the rest of TIA.  There is probably a 
--                lot of stuff that can be eliminated later.  Also,
--                keep in mind that some of this is not good when doing
--                high speed design!
--
--   !!!!!!!!!!! CLEAN THIS CODE UP PRIOR TO RELEASE!!!!  !!!!!!!!!!!!!!!!!!
--
--   Date      :  January 12, 2005
--                
-------------------------------------------------------------------------------

library IEEE;
    use IEEE.std_logic_1164.all;
    use IEEE.std_logic_unsigned.all;
    use IEEE.std_logic_arith.all;

library A2600;
    use A2600.tia_pkg.all;
    -- synthesis translate_off
    use A2600.tia_sim_comps.all;
    -- synthesis translate_on

entity tia_ctl_pf is
port
(

   -- Clock and system reset 
   clk          : in  std_logic; -- Main system clock 
   reset_sys    : in  std_logic; -- Primary reset

   -- Reference enable inputs to sync
   -- system clock to actual TIA rates.
   ena_sys      : in  std_logic;
   ena_pix      : in  std_logic;

   -- Simulation only reference signals
   -- synthesis translate_off
   ref_sys_clk  : in  std_logic;
   ref_pix_clk  : in  std_logic;
   ref_newline  : out std_logic;
   -- synthesis translate_on
   
   -- RSYNC strobe from regfile
   rsync        : in  std_logic;

   -- WSYNC strobe from regfile
   wsync        : in  std_logic;

   -- VSYNC & VBLANK register inputs from regfile
   vsync        : in  std_logic;
   vblank       : in  std_logic;

   -- Horizontal move strobe from regfile
   hmove        : in  std_logic;

   -- Playfield register inputs
   pf0          : in  std_logic_vector(3 downto 0);
   pf1          : in  std_logic_vector(7 downto 0);
   pf2          : in  std_logic_vector(7 downto 0);

   -- Playfield reflect bit from regfile
   pf_ref       : in  std_logic;

   -- Horizontal motion input vectors
   hmp0         : in  std_logic_vector(3 downto 0);
   hmp1         : in  std_logic_vector(3 downto 0);
   hmm0         : in  std_logic_vector(3 downto 0);
   hmm1         : in  std_logic_vector(3 downto 0);
   hmbl         : in  std_logic_vector(3 downto 0);

   -- CPU clock reference
   cpu_clk      : in  std_logic;

   -- CPU clock reset control
   ctl_rst_cpu  : out std_logic;

   -- CPU ready signal 
   cpu_rdy      : out std_logic;

   -- Playfield graphics output
   pf_out       : out std_logic;

   -- Playfield Center Delayed
   cntd         : out std_logic;

   -- Signals driven to video control logic
   vid_csync    : out std_logic;
   vid_hsync    : out std_logic;
   vid_vsync    : out std_logic;
   vid_cburst   : out std_logic;
   vid_blank    : out std_logic;
   vid_hblank   : out std_logic;

   -- The following signals are related to horizontal
   -- motion.  These are to be used as simulation
   -- references in the event something goes wrong...
   -- synthesis translate_off
   ref_motclk   : out std_logic;
   ref_en_blm_n : out std_logic;
   ref_en_p0m_n : out std_logic;
   ref_en_m0m_n : out std_logic;
   ref_en_p1m_n : out std_logic;
   ref_en_m1m_n : out std_logic;
   -- synthesis translate_on

   -- This signal allows the object counters
   -- to advance (i.e. draw the things!)
   adv_obj      : out std_logic;

   -- These are the motion signals used
   -- in the synthesizable application...see
   -- objects for details.
   ball_mot     : out std_logic;
   p0_mot       : out std_logic;
   m0_mot       : out std_logic;
   p1_mot       : out std_logic;
   m1_mot       : out std_logic;

   -- Finally, the audio clock signals
   aud_clk1     : out std_logic;
   aud_clk2     : out std_logic 

);
end tia_ctl_pf;

architecture rtl of tia_ctl_pf is

   -- The time that H1 and H2 would fire are indicated
   -- by these signals.
   signal h1_clk            : std_logic;
   signal h2_clk            : std_logic;

   -- Internal flop enable signals
   signal h1_ena            : std_logic;
   signal h2_ena            : std_logic;

   -- Current sequencing count
   signal cur_cnt           : seq_int; 

   -- Control signals generated by the horizontal timing
   -- sequence counter.
   signal shs_i             : std_logic;
   signal rhs_i             : std_logic;
   signal rcb_i             : std_logic;
   signal rhb_i             : std_logic;
   signal lrhb_i            : std_logic;
   signal cnt_i             : std_logic;
   signal end_i             : std_logic;

   -- The set hblank flop that also
   -- resets the sequence counter.
   signal shb               : std_logic;

   -- Output of RSYNC RS latch
   signal rsyn_lat          : std_logic;

   -- Input to the rsync flip flop
   signal rsync_input       : std_logic;

   -- CPU clock sync signal (sync'ed to H1 clock).
   signal rsynd             : std_logic;

   -- Internal resets
   signal reset_sequencer   : std_logic;
   signal reset_seqclk      : std_logic;
   signal reset_synclat     : std_logic;

   -- Internal registers (i.e. register output)
   signal rst_hs            : std_logic; -- Reset hsync
   signal hsync_r           : std_logic; -- Horizontal sync reg
   signal rcb               : std_logic; -- Color burst delayed reg
   signal blank             : std_logic; -- Common blank signal

   -- Ready latch signals
   signal rdy_lat_set       : std_logic;
   signal rdy_lat_clr       : std_logic;
   signal rdy_n             : std_logic;

   -- Signals involved in horizontal movement
   signal sec_lat_out         : std_logic; -- output of SEC latch
   signal hmove_dcnt          : std_logic_vector(3 downto 0); -- Hmove ref. cnt
   signal en_dcnt             : std_logic; -- downcount enable
   signal nx1, nx2, nx3       : std_logic; -- nodes in 3 NMOS latch chain
   signal nx1_c, nx2_c, nx3_c : std_logic; -- nodes in 3 NMOS latch chain
   signal nx1_s, nx2_s, nx3_s : std_logic; -- nodes in 3 NMOS latch chain
   signal sec                 : std_logic; -- SEC pulse
   signal reset_seclat        : std_logic; -- clears SEC latch

   -- Audio clock pre-flop references...
   signal aud_clk1_i        : std_logic;
   signal aud_clk2_i        : std_logic;

   -- The "invert MSB" motion values for 
   -- the motion comparitors...
   signal cmp_hmp0          : std_logic_vector(3 downto 0);
   signal cmp_hmp1          : std_logic_vector(3 downto 0);
   signal cmp_hmm0          : std_logic_vector(3 downto 0);
   signal cmp_hmm1          : std_logic_vector(3 downto 0);
   signal cmp_hmbl          : std_logic_vector(3 downto 0);

   -- Stop motion signals!
   signal stopm_p0          : std_logic;
   signal stopm_p1          : std_logic;
   signal stopm_m0          : std_logic;
   signal stopm_m1          : std_logic;
   signal stopm_bl          : std_logic;

   -- Internal motion enable bits...
   signal mot_ena_p0        : std_logic;
   signal mot_ena_p1        : std_logic;
   signal mot_ena_m0        : std_logic;
   signal mot_ena_m1        : std_logic;
   signal mot_ena_bl        : std_logic;

   -- Signals used to generate the HBLANK signal
   signal clr_hblank_lat    : std_logic; -- Clears the HBLANK latch
   signal clr_hblank_lat_normal    : std_logic;
   signal regular_hblank    : std_logic; -- "hblank fires normally"
   signal late_hblank       : std_logic; -- "hblank fires 8 cycles late"
   signal gate_regular      : std_logic; -- AND gate indicating reg. blank
   signal gate_late         : std_logic; -- AND gate indicating late blank
   signal hblank_i          : std_logic; -- internal horiz. blank signal
   signal reset_hbl_flop    : std_logic; -- clears the HBLANK flop
   signal hblank_n          : std_logic; -- output of HBLANK flop!

   -- Signals dealing with playfield serialization
   signal playfield         : std_logic_vector(19 downto 0);
   signal up_shift          : std_logic_vector(19 downto 0);
   signal down_shift        : std_logic_vector(19 downto 0);
   signal pf_up             : std_logic;
   signal pf_down           : std_logic;
   signal pf_up_out         : std_logic;
   signal pf_down_out       : std_logic;

   -- synthesis translate_off
   -- Silly reference signals...none are synthsized...
   -- use these to compare "expected" against "real"
   signal ref_pix_cnt       : integer;
   -- synthesis translate_on

begin

   ------------------------------------------------------
   -- This component generates all our silly sequencing
   -- logic for this circuit...
   ------------------------------------------------------
   horiz_seq_0 : tia_sequencer
   port map
   (

      -- synthesis translate_off
      sim_clk   => ref_sys_clk,
      -- synthesis translate_on
      clk       => clk,
      reset_sys => reset_sys,
      enable    => ena_sys,
      reset_ctr => reset_sequencer,
      rlat_in   => reset_seqclk,
      p1_clk    => h1_clk,
      p2_clk    => h2_clk,
      p1_ena    => h1_ena,
      p2_ena    => h2_ena,
      cnt_out   => cur_cnt,
      rlat_out  => rsyn_lat,
      tap_out   => open

   );

   ------------------------------------------------------
   -- This gate generates the reset for the CPU clock
   -- Be aware that h2_clk is not a clock in the "FPGA"
   -- sense...it is actually the output of a counter!
   ------------------------------------------------------
   ctl_rst_cpu <= (rsynd and h2_clk);

   -------------------------------------------------------
   -- SHB clears the sequence counter...the sequence
   -- counter requires a funky pseudo-asynchronous reset.
   -- See the sequencer logic for details.
   -------------------------------------------------------
   reset_sequencer <= shb;

   -----------------------------------------------------------------------
   -- This gate resets the sequencer clocking.  It also appears
   -- to play a role in sync'ing the sequencer to the CPU clock :
   -- 
   --                              This is RSYNC tied to NMOS pulldown.
   --                              If the CPU clock is high, then the
   --                              pulldown yanks rsync to ground. 
   -----------------------------------------------------------------------
   reset_seqclk    <= reset_sys or (rsync and not(cpu_clk));

   ------------------------------------------------------
   -- This process asserts control signals depending on
   -- the state of the seq_cnt process above.  Note that
   -- this process creates combinational logic...
   ------------------------------------------------------
   process(cur_cnt)
   begin

       -- By default, keep these guys off...
       shs_i  <= '0';
       rhs_i  <= '0';
       rcb_i  <= '0';
       rhb_i  <= '0';
       lrhb_i <= '0';
       cnt_i  <= '0';
       end_i  <= '0';

       -- Decode the output of the sequence counter so that we 
       -- can properly assert various control signals.
       case cur_cnt is

            when  SET_HSYNC_CNT     => shs_i  <= '1';
            when  RESET_HSYNC_CNT   => rhs_i  <= '1';
            when  COLORBURST_CNT    => rcb_i  <= '1';
            when  RESET_HBLANK      => rhb_i  <= '1';
            when  LATE_RESET_HBLANK => lrhb_i <= '1';
            when  CENTER_CNT        => cnt_i  <= '1';
            when  END_SEQ_CNT       => end_i  <= '1';

            -- Default case sets all control signals low.
            when  OTHERS            => shs_i  <= '0';
                                       rhs_i  <= '0';
                                       rcb_i  <= '0';
                                       rhb_i  <= '0';
                                       lrhb_i <= '0';
                                       cnt_i  <= '0';
                                       end_i  <= '0';
       end case;

   end process;

   ----------------------------------------------------
   -- It appears that we need a funky construct to
   -- properly emulate the nice rsynd / shb latch.
   -- If we only needed to reset the sequencer upon
   -- a receipt of end_i, then we'd have no problem
   -- emulating the latch with edge-triggered devices 
   -- w. enable since that signal is sync'ed to H2.
   --
   -- Unfortunately, as with everything in TIA, we
   -- need to do something a little more clever.
   -- rsyn_lat can arrive at a bunch of silly different
   -- times causing the universe to end in some cases.
   --
   -- We need to have both a combinational and 
   -- sequential component to latch this as seen
   -- below...the timing of a counter reset appears to
   -- be very critical (i.e. I had lots of filthy bugs 
   -- when clearing counters)!
   --
   -- By the way, this is when I decided to make the
   -- nutty little "tia_d_flop" component.
   ----------------------------------------------------

   -- Create reset
   rsync_input <= end_i or rsyn_lat;

   -- Dual phase flop to drive RSYN related signals
   rsync_flop : tia_d_flop
   generic map(
      flop_style => REGULAR_D
   )
   port map
   (

      clk          => clk,
      reset        => reset_sys,
      reset_gate   => '0',
      p1_clk       => h1_clk,
      p2_clk       => h2_clk,
      data_in      => rsync_input,

      -- D-Flop outputs based on phase
      p1_out       => rsynd,
      p2_out       => shb

   );

   ----------------------------------------------
   -- Various signals that require an H2 phase
   -- delay....these are reset by the "power on"
   -- reset signal...nothing else in TIA clears 
   -- them out!
   ----------------------------------------------

   -- Instantiate the flop for center delayed
   cntd_flop : tia_d_flop
   generic map(
      flop_style => REGULAR_D
   )
   port map
   (

      clk          => clk,
      reset        => reset_sys,
      reset_gate   => '0',
      p1_clk       => h1_clk,
      p2_clk       => h2_clk,
      data_in      => cnt_i,

      -- D-Flop outputs based on phase
      p1_out       => open,
      p2_out       => cntd -- Center Delayed

   );

   reset_hsync_flop : tia_d_flop
   generic map(
      flop_style => REGULAR_D
   )
   port map
   (

      clk          => clk,
      reset        => reset_sys,
      reset_gate   => '0',
      p1_clk       => h1_clk,
      p2_clk       => h2_clk,
      data_in      => rhs_i,

      -- D-Flop outputs based on phase
      p1_out       => open,
      p2_out       => rst_hs -- Reset hsync flop

   );

   -- Generate the or gates for audio clock generation
   aud_clk1_i <= rhs_i  or cnt_i;
   aud_clk2_i <= lrhb_i or shb;

   -- Instantiate audio clock flops
   aud1_flop : tia_d_flop
   generic map(
      flop_style => REGULAR_D
   )
   port map
   (

      clk          => clk,
      reset        => reset_sys,
      reset_gate   => '0',
      p1_clk       => h1_clk,
      p2_clk       => h2_clk,
      data_in      => aud_clk1_i,

      -- D-Flop outputs based on phase
      p1_out       => open,
      p2_out       => aud_clk1 -- Audio clock 1 reference

   );

   aud2_flop : tia_d_flop
   generic map(
      flop_style => REGULAR_D
   )
   port map
   (

      clk          => clk,
      reset        => reset_sys,
      reset_gate   => '0',
      p1_clk       => h1_clk,
      p2_clk       => h2_clk,
      data_in      => aud_clk2_i,

      -- D-Flop outputs based on phase
      p1_out       => open,
      p2_out       => aud_clk2 -- Audio clock 2 reference

   );

   ----------------------------------------------------------
   -- These components register other single cycle (H2) delay
   -- signals.  The difference here is that other signals
   -- reset these flip flops...
   ----------------------------------------------------------

   -- First, create the reset
   reset_synclat <= rst_hs or reset_sys;

   -- Instantiate the flop for colorburst
   colorb_flop : tia_d_flop
   generic map(
      flop_style => FEEDBK_RST
   )
   port map
   (

      clk          => clk,
      reset        => reset_sys,
      reset_gate   => reset_synclat,
      p1_clk       => h1_clk,
      p2_clk       => h2_clk,
      data_in      => rcb_i,

      -- D-Flop outputs based on phase
      p1_out       => open,
      p2_out       => rcb

   );

   -- Instantiate the flop for hsync
   hsync_flop : tia_d_flop
   generic map(
      flop_style => FEEDBK_RST
   )
   port map
   (

      clk          => clk,
      reset        => reset_sys,
      reset_gate   => reset_synclat,
      p1_clk       => h1_clk,
      p2_clk       => h2_clk,
      data_in      => shs_i,

      -- D-Flop outputs based on phase
      p1_out       => open,
      p2_out       => hsync_r

   );

   --------------------------------
   -- Playfield generation logic --
   --------------------------------

   -- Here we do a simple remapping of the playfield bits
   -- so that the "normal" and "reflected" outputs are a 
   -- little easier to manage!
   playfield(0)  <= pf0(0); -- PF0 4
   playfield(1)  <= pf0(1); -- PF0 5
   playfield(2)  <= pf0(2); -- PF0 6
   playfield(3)  <= pf0(3); -- PF0 7
   playfield(4)  <= pf1(7); -- PF1 7
   playfield(5)  <= pf1(6); -- PF1 6
   playfield(6)  <= pf1(5); -- PF1 5
   playfield(7)  <= pf1(4); -- PF1 4
   playfield(8)  <= pf1(3); -- PF1 3
   playfield(9)  <= pf1(2); -- PF1 2
   playfield(10) <= pf1(1); -- PF1 1
   playfield(11) <= pf1(0); -- PF1 0
   playfield(12) <= pf2(0); -- PF2 0
   playfield(13) <= pf2(1); -- PF2 1
   playfield(14) <= pf2(2); -- PF2 2
   playfield(15) <= pf2(3); -- PF2 3
   playfield(16) <= pf2(4); -- PF2 4
   playfield(17) <= pf2(5); -- PF2 5
   playfield(18) <= pf2(6); -- PF2 6
   playfield(19) <= pf2(7); -- PF2 7
   
   -- This process shifts playfield data out of the playfield
   -- registers.  The playfield registers seem to be clocked
   -- out using a type of "token".  This token is dropped into
   -- the registers @ the time rhb_i is asserted as well as the
   -- time cnt_i is asserted.  The reflection bit determines the
   -- direction to clock data out when cnt_i is asserted.  Data
   -- is always output normally when rhb_i is asserted.

   -- Yes, we could probably implement this with a simple counter
   -- that muxes out data (this would probably save area too), but 
   -- that's no fun!

   -- First generate the up/down enable signals
   pf_up   <= rhb_i or (cnt_i and not(pf_ref)); -- Don't reflect.
   pf_down <= pf_ref and cnt_i;                 -- Reflect playfield if true.

   -- Process for the shift registers / serialization of playfield
   process(clk, reset_sys)
   begin

       if (reset_sys = '1') then

           up_shift    <= (others => '0');
           down_shift  <= (others => '0');
           pf_up_out   <= '0';
           pf_down_out <= '0';

       elsif(clk'event and clk = '1') then

           -- Prepare to determine the bit present on the 
           -- H@ phase of the clock;
           if (h2_ena = '1') and (ena_sys = '1') then

               -- Always shift the enable bit into the appropriate
               -- shift register...
               up_shift(1)    <= pf_up;
               down_shift(18) <= pf_down;

               -- This logic controls "normal" playfield serialization
               if (pf_up = '1') then

                   pf_up_out <= playfield(0);

               else

                   -- By default, drive a zero out...
                   pf_up_out    <= '0';

                   -- Here we see what the value of the playfield
                   -- bit should be in the playfield serial stream.
                   for i in 1 to 19 loop

                      -- See if we should drive a '1' out in the 
                      -- playfield serial stream.
                      if ((up_shift(i) and playfield(i)) = '1') then
                         pf_up_out <= '1';
                      end if;

                      -- Shift the bit to the next enable
                      up_shift(i)   <= up_shift(i-1);

                   end loop;

                   -- To keep warnings from being generated, 
                   -- clear out up_shift(0)
                   up_shift(0) <= '0';

               end if;

               -- Reflected playfield serialization logic...
               if (pf_down = '1') then
                      
                   pf_down_out <= playfield(19);

               else

                   -- By default, drive a zero out...
                   pf_down_out    <= '0';

                   -- Here we see what the value of the playfield
                   -- bit should be in the playfield serial stream.
                   for i in 18 downto 0 loop

                      -- See if we should drive a '1' out in the 
                      -- playfield serial stream.
                      if ((down_shift(i) and playfield(i)) = '1') then
                         pf_down_out <= '1';
                      end if;

                      -- Shift the bit to the next enable
                      down_shift(i)   <= down_shift(i+1);

                   end loop;
                      
                   -- To keep warnings from being generated, 
                   -- clear out down_shift(19)
                   down_shift(19) <= '0';

               end if;

           end if;

       end if;

   end process;

   -- Process to clock out serialized playfield data...
   -- This should be register delay matched to hblank.
   -- Use ref_pix_cnt to verify.
   process(clk, reset_sys)
   begin

         if (reset_sys = '1') then
             pf_out <= '0';
         elsif(clk'event and clk = '1') then
             if (ena_pix = '1') then
                pf_out <= pf_up_out or pf_down_out;
             end if;
         end if;

   end process;

   ---------------------------------------------------------------
   -- The following processes are the horizontal motion control
   -- processes!  These drive extra clock cycles to the object
   -- counters so that objects move under hardware assist.  We 
   -- must also preserve a bug in this logic that continues to 
   -- stuff extra cycles creating the "Cosmic Ark" starfield 
   -- effect...we'll discuss that later...
   ---------------------------------------------------------------
   
   -- First, we need a latch that is responsible for creating the
   -- SEC pulse upon assertion of the HMOVE signal...
   hmove_latch_0 : tia_latch
   port map(

        clk    => clk,
        set    => hmove,
        clear  => reset_seclat,
        output => sec_lat_out
   );

   -- The following needs to be implemented in the fine
   -- TIA half sequential / half combinational style...

   -- By the way, clear the latch any time nx3 is high or
   -- when a system reset is present...
   reset_seclat <= nx3 or reset_sys;

   -- Now the SEC pulse generator...
   
   -- Combinational component for SEC generation
   process(sec_lat_out, nx1, nx2)
   begin

       nx1_c <= not(sec_lat_out);
       nx2_c <= not(nx1);
       nx3_c <= nx2;

   end process;

   -- Sequential component for SEC generation
   process(clk, reset_sys)
   begin

      if (reset_sys = '1') then

          nx1_s <= '1';
          nx2_s <= '0';
          nx3_s <= '0';

      elsif(clk'event and clk = '1') then

          -- Clocked on H1 phase
          if (h1_clk = '1') then
             nx1_s <= nx1_c;
             nx3_s <= nx3_c;
          end if;

          -- Clocked on H2 phase
          if (h2_clk = '1') then
            nx2_s <= nx2_c;
          end if;

      end if;

   end process;

   -- Generate pulse signals here...
   nx1 <= nx1_c when (h1_clk = '1') else nx1_s;
   nx2 <= nx2_c when (h2_clk = '1') else nx2_s;
   nx3 <= nx3_c when (h1_clk = '1') else nx3_s;
   
   -- The SEC signal is simply nx2.
   sec <= nx2;

   -- Next, we need a reference counter.  This downcounter
   -- is triggered by SEC, counts to zero, and then waits for the
   -- next SEC pulse to arrive!  It downcounts on each H2 phase 
   -- of the clock.
   process(clk, reset_sys)
   begin

       if (reset_sys = '1') then

           hmove_dcnt <= "1111";
           en_dcnt    <= '0';

       elsif (clk'event and clk = '1') then

           -- When H2 is present....
           if (h2_ena = '1') and (ena_sys = '1') then

               -- Any time we see SEC or the downcount enable
               -- asserted, decrement the counter...
               if (sec = '1') or (en_dcnt = '1') then

                   en_dcnt <= '1';
                   hmove_dcnt <= hmove_dcnt - 1;

               end if;

               -- Once we see the counter at zero, reset
               -- the counter and clear the enable downcount 
               -- flag!
               if (hmove_dcnt = "0000") then

                   hmove_dcnt <= "1111";
                   en_dcnt    <= '0';

               end if;

           end if;

       end if;

   end process;

   -- Let's generate the logic that will stop horizontal motion
   -- based on the value the program dictates...

   -- Here we invert the MSB of the motion values latched in
   -- the write register logic.
   process(hmp0, hmp1, hmm0, hmm1, hmbl)
   begin
       cmp_hmp0 <= not(hmp0(3)) & hmp0(2 downto 0);
       cmp_hmp1 <= not(hmp1(3)) & hmp1(2 downto 0);
       cmp_hmm0 <= not(hmm0(3)) & hmm0(2 downto 0);
       cmp_hmm1 <= not(hmm1(3)) & hmm1(2 downto 0);
       cmp_hmbl <= not(hmbl(3)) & hmbl(2 downto 0);
   end process;

   -- Now generate the signals that stop the object advance
   -- latches...this is a combinational circuit!
   process(hmove_dcnt, cmp_hmp0, cmp_hmp1, cmp_hmm0, cmp_hmm1, cmp_hmbl)
   begin

       -- Stop player 0 motion
       if (cmp_hmp0 /= not(hmove_dcnt)) then
          stopm_p0 <= '0';
       else
          stopm_p0 <= '1';
       end if;

       -- Stop player 1 motion
       if (cmp_hmp1 /= not(hmove_dcnt)) then
          stopm_p1 <= '0';
       else
          stopm_p1 <= '1';
       end if;

       -- Stop missile 0 motion
       if (cmp_hmm0 /= not(hmove_dcnt)) then
          stopm_m0 <= '0';
       else
          stopm_m0 <= '1';
       end if;

       -- Stop missile 1 motion
       if (cmp_hmm1 /= not(hmove_dcnt)) then
          stopm_m1 <= '0';
       else
          stopm_m1 <= '1';
       end if;

       -- Stop...heh..heh...ball motion...heh...heh
       if (cmp_hmbl /= not(hmove_dcnt)) then
          stopm_bl <= '0';
       else
          stopm_bl <= '1';
       end if;

   end process;

   -- With all the above in place, we can generate the motion
   -- enable signals...
   process(clk, reset_sys)
   begin

        if (reset_sys = '1') then

            mot_ena_p0 <= '0';
            mot_ena_p1 <= '0';
            mot_ena_m0 <= '0';
            mot_ena_m1 <= '0';
            mot_ena_bl <= '0';

        elsif(clk'event and clk = '1') then

            if (ena_sys = '1') then 

               -- Set the enables for the silly
               -- motion enable signal when necessary...
               if (sec = '1') and (h1_clk = '1') then

                   mot_ena_p0 <= '1';
                   mot_ena_p1 <= '1';
                   mot_ena_m0 <= '1';
                   mot_ena_m1 <= '1';
                   mot_ena_bl <= '1';

               end if;

               -- Clear the motion enable signals
               -- when necessary...this is done when the
               -- H1 clock is active...

               -- Player 0
               if (h1_clk = '1') and (stopm_p0 = '1') then
                  mot_ena_p0 <= '0';
               end if;

               -- Player 1
               if (h1_clk = '1') and (stopm_p1 = '1') then
                  mot_ena_p1 <= '0';
               end if;

               -- Missile 0
               if (h1_clk = '1') and (stopm_m0 = '1') then
                  mot_ena_m0 <= '0';
               end if;
 
               -- Missile 1
               if (h1_clk = '1') and (stopm_m1 = '1') then
                  mot_ena_m1 <= '0';
               end if;

               -- Heh heh ... Ball
               if (h1_clk = '1') and (stopm_bl = '1') then
                  mot_ena_bl <= '0';
               end if;
  
            end if;

        end if;

   end process;

   -- Output clock enable signals for the objects...
   adv_obj  <= hblank_n;
   ball_mot <= mot_ena_bl and h1_ena;
   p0_mot   <= mot_ena_p0 and h1_ena;
   m0_mot   <= mot_ena_m0 and h1_ena;
   p1_mot   <= mot_ena_p1 and h1_ena;
   m1_mot   <= mot_ena_m1 and h1_ena;
   
   ---------------------------------------------------------------
   -- The following logic generates the horizontal blank signal --
   ---------------------------------------------------------------
   
   -- First, this latch is set by "set hblank" and cleared
   -- by the SEC pulse.  It appears that if the SEC pulse
   -- clears this latch, hblank is not set until "late
   -- reset hblank" arrives (i.e. motion).

   clr_hblank_lat <= sec or reset_sys;
   clr_hblank_lat_normal <= rhb_i or reset_sys;

   hblank_latch_0 : tia_latch
   port map(

        clk    => clk,
        set    => shb,
        clear  => clr_hblank_lat,
        output => regular_hblank -- normal hblank if high
   );

   hblank_latch_1 : tia_latch
   port map(

        clk    => clk,
        set    => shb,
        clear  => clr_hblank_lat_normal,
        output => vid_hblank -- normal hblank if high
   );

   -- This indicates that we fire hblank late
   late_hblank  <= not(regular_hblank);

   -- Now that we know which blank to pay attention to, create
   -- the gates that shall drive the hblank sequential logic!
   gate_regular <= rhb_i        and regular_hblank;
   gate_late    <= lrhb_i       and late_hblank;
   hblank_i     <= gate_regular or  gate_late;

   -- Next is the hblank flip-flop...

   -- This generates the reset for this flop...
   reset_hbl_flop <= reset_sys or shb;   

   -- This is the flip flop (i.e. nor based with feedback loop)
   -- that stores the current hblank value.
   hblank_flop : tia_d_flop
   generic map(
      flop_style => FEEDBK_RST
   )
   port map
   (

      clk          => clk,
      reset        => reset_sys,
      reset_gate   => reset_hbl_flop,
      p1_clk       => h1_clk,
      p2_clk       => h2_clk,
      data_in      => hblank_i,

      -- D-Flop outputs based on phase
      p1_out       => open,
      p2_out       => hblank_n

   );
   
   ---------------------------------------------------------------
   -- This latch generates the CPU ready signal.  This latch is
   -- used to keep the CPU in sync with the TIA.  First we need
   -- to generate the control signals.... 
   ---------------------------------------------------------------

   -- The latch is cleared when the input clock (inverted) and
   -- set horizontal blank are true...the reference signal for
   -- the system clock is the same as the "actual" system clock
   -- inverted...
   rdy_lat_clr <= (ena_sys and shb) or reset_sys;

   -- The latch is set when the WSYNC strobe is present and
   -- the set horizontal blank signal is not asserted.  My guess
   -- is that this gate was necessary to prevent a race condition.
   -- Actually, this is to prevent a wait state if the counter
   -- is at the first count of the line....why waste a whole line?
   rdy_lat_set <= not(shb) and wsync;

   -- And now, the latch...
   rdy_latch_0 : tia_latch
   port map(

        clk    => clk,
        set    => rdy_lat_set,
        clear  => rdy_lat_clr,
        output => rdy_n
   );

   -- And, finally, invert the output of the latch.
   cpu_rdy <= not(rdy_n);

   -- This process registers the blank signal on the pixel clock
   process(clk, reset_sys)
   begin

       if (reset_sys = '1') then
           blank <= '0';
       elsif(clk'event and clk = '1') then
           if (ena_pix = '1') then
               blank <= not(hblank_n) or vblank;
           end if;
       end if;

   end process;

   --------------------------------------------------------------
   -- Here we generate all those signals going to the video
   -- control logic.  Yes, some signals are being replicated,
   -- but this is done basically for readibility.  Some of these
   -- are quite possibly useless...I left them all here just
   -- in case someone wants to use them!
   --------------------------------------------------------------
   vid_csync    <= hsync_r xnor vsync; -- Composite sync
   vid_hsync    <= hsync_r;            -- Horizontal sync
   vid_vsync    <= vsync;              -- Vertical sync
   vid_cburst   <= vsync   nor rcb;    -- Colorburst (probably uesless)
   vid_blank    <= blank;              -- Gated & registered blank signal
    
   -----------------------------------------------------
   --                                                 --
   --      END OF CODE TARGETED FOR SYNTHESIS!!!!     --
   --                                                 --
   -----------------------------------------------------

   -----------------------------------------------------------
   -- Sleek, silly, simulation reference....none of this is 
   -- to be synthesized...these are used to insure timing is
   -- correct with respect to the H1 and H2 reference clocks.
   -----------------------------------------------------------

   -- synthesis translate_off

   -- Newline reference for testing purposes
   ref_newline <= shb;

   -- Count the cycles where blank is not active to see if it
   -- equals 160...this would also be useful for debugging games
   process(ref_pix_clk, reset_sys, blank)
   begin

       if (reset_sys = '1') or (blank = '1') then
           ref_pix_cnt <= 0;
       elsif(ref_pix_clk'event and ref_pix_clk = '1') then

           if (blank = '0') then
               ref_pix_cnt <= ref_pix_cnt + 1;
           end if;

       end if;

   end process;

   -- Generate the motion clock...for reference
   ref_motclk <= not(hblank_n) nor ref_sys_clk; -- Clock gating is bad...that's
                                                -- why this is not synthesized. This
                                                -- is how TIA generates the clock.

   -- This component simulates the horizontal motion logic
   -- at the gate level. I left this in here since it's
   -- tons of fun to mimic perfectly.
   --hmotion_sim_0 : tia_hmotion_sim
   --port map
   --(

   --   h1_clk     => h1_clk,
   --   h2_clk     => h2_clk,
   --   reset      => reset_sys,

   --   hmove      => hmove,

   --   p0_vec     => hmp0,
   --   p1_vec     => hmp1,
   --   m0_vec     => hmm0,
   --   m1_vec     => hmm1,
   --   bl_vec     => hmbl,


   --   p0_ec_n    => ref_en_p0m_n,
   --   p1_ec_n    => ref_en_p1m_n,
   --   m0_ec_n    => ref_en_m0m_n,
   --   m1_ec_n    => ref_en_m1m_n,
   --   bl_ec_n    => ref_en_blm_n 

   --);

   -- synthesis translate_on

end rtl;
