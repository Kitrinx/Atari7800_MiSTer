`define CS_NONE     'h0
`define CS_RAM0     'h1
`define CS_RAM1     'h2
`define CS_RIOT_IO  'h3
`define CS_RIOT_RAM 'h4
`define CS_TIA      'h5
`define CS_BIOS     'h6
`define CS_MARIA    'h7
`define CS_CART     'h8

`define chipselect  logic[3:0]

//`define SIM