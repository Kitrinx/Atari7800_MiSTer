`timescale 1ns / 1ps

module audio(input logic [3:0] AUDC0, AUDC1,
	         input logic [4:0] AUDF0, AUDF1,
	         input logic CLK_30, //30khz clock
	         output logic AUD0,AUD1
	         );

	logic [4:0] counter0, counter1 = 5'b0;
	integer rep0,rep1,ind0,ind1 = 0;
	logic [1:0] pattern45 = 2'b10;
	logic pattern0b = 1'b1;
	logic [14:0] pattern1 = 15'b111100010011010;
	logic [30:0] pattern6a = 31'b1111111111111111110000000000000;
	logic [30:0] pattern79 = 31'b1111100011011101010000100101100;
	logic [5:0] patterncd = 6'b111000;
	logic [92:0] patterne =  93'b111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000;
	logic [92:0] patternf =  93'b111111111100000111000000011110000000000111111000111111000011111111100000011111000000111100000;
	logic [464:0] pattern2 = 465'b111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000001111111111111111111111111111111000000000000000000111111111111100000000000000000011111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000111111111111111111111111111111100000000000001111111111111111110000000000000;
	logic [464:0] pattern3 = 465'b111111000000100011100111110001111111000111100011001100000111111111000100000111011001111111111100000100000111010011111111111100000100111110010111111111111000000100111110110111111111100000011100110000100111111000000000010000110111101111110000000000110000110100001111100000000011100011110101111111100000111110000011110101111111100001100000000111000101111111000011000000011111011101111111000010000111111110010001111000000010001111111000110111111000000110011110000011100;
	logic [510:0] pattern8 = 511'b1111111110000011110111110001011100110010000010010100111011010001111001111100110110001010100100011100011011010101110001001100010001000000001000010001100001001110010101011000011011110100110111001000101000010101101001111110110010010010110111111001001101010011001100000001100011001010001101001011111110100010110001110101100101100111100011111011101000001101011011011101100000101101011111010101010000001010010101111001011101110000001110011101001001111010111010100010010000110011100001011110110110011010000111011110000;

	always_comb begin
		case (AUDC0)
			4'h0,4'hb: rep0 = 1;
			4'h1: rep0 = 15;
			4'h2,4'h3: rep0 = 465;
			4'h4,4'h5: rep0 = 2;
			4'h6,4'h7,4'h9,4'ha: rep0 = 31;
			4'h8: rep0 = 511;
			4'hc,4'hd: rep0 = 6;
			4'he,4'hf: rep0 = 93;
			default: rep0 = 1;
		endcase
		case (AUDC1)
			4'h0,4'hb: rep1 = 1;
			4'h1: rep1 = 15;
			4'h2,4'h3: rep1 = 465;
			4'h4,4'h5: rep1 = 2;
			4'h6,4'h7,4'h9,4'ha: rep1 = 31;
			4'h8: rep1 = 511;
			4'hc,4'hd: rep1 = 6;
			4'he,4'hf: rep1 = 93;
			default: rep0 = 1;
		endcase
	end

	always_ff @(posedge CLK_30) begin //divide the clk by the frequency value
		if (counter0 == AUDF0) begin
			case (AUDC0)
                    4'h0,4'hb: AUD0 <= pattern0b;
                    4'h1: AUD0 <= pattern1[ind0];
                    4'h2: AUD0 <= pattern2[ind0];
                    4'h3: AUD0 <= pattern3[ind0];
                    4'h4,4'h5: AUD0 <= pattern45[ind0];
                    4'h6,4'ha: AUD0 <= pattern6a[ind0];
                    4'h7,4'h9: AUD0 <= pattern79[ind0];
                    4'h8: AUD0 <= pattern8[ind0];
                    4'hc,4'hd: AUD0 <= patterncd[ind0];
                    4'he: AUD0 <= patterne[ind0];
                     4'hf: AUD0 <= patternf[ind0];
                     default: AUD0 <= 1'bx;
                 endcase
            ind0 <= (ind0 + 1) % rep0;
			counter0 <= 0;
		end
		else
			counter0 <= counter0 + 1'd1;

		if (counter1 == AUDF1) begin
			case (AUDC1)
                    4'h0,4'hb: AUD1 <= pattern0b;
                    4'h1: AUD1 <= pattern1[ind1];
                    4'h2: AUD1 <= pattern2[ind1];
                    4'h3: AUD1 <= pattern3[ind1];
                    4'h4,4'h5: AUD1 <= pattern45[ind1];
                    4'h6,4'ha: AUD1 <= pattern6a[ind1];
                    4'h7,4'h9: AUD1 <= pattern79[ind1];
                    4'h8: AUD1 <= pattern8[ind1];
                    4'hc,4'hd: AUD1 <= patterncd[ind1];
                    4'he: AUD1 <= patterne[ind1];
                     4'hf: AUD1 <= patternf[ind1];
                     default: AUD1 <= 1'bx;
                 endcase
            ind1 <= (ind1 + 1) % rep1;
			counter1 <= 0;
		end
		else
			counter1 <= counter1 + 1'd1;
	end


endmodule:  audio
